library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all; 

entity chippy_bcd_lut is
	port (addr : in std_logic_vector(7 downto 0);
		data : out std_logic_vector(11 downto 0) );
end chippy_bcd_lut;		   

architecture behavioural of chippy_bcd_lut is
begin
	process(addr)
	begin
		if addr = 0 then data <="000000000000";
		elsif addr = 1 then data <="000000000001";
		elsif addr = 2 then data <="000000000010";
		elsif addr = 3 then data <="000000000011";
		elsif addr = 4 then data <="000000000100";
		elsif addr = 5 then data <="000000000101";
		elsif addr = 6 then data <="000000000110";
		elsif addr = 7 then data <="000000000111";
		elsif addr = 8 then data <="000000001000";
		elsif addr = 9 then data <="000000001001";
		elsif addr = 10 then data <="000000010000";
		elsif addr = 11 then data <="000000010001";
		elsif addr = 12 then data <="000000010010";
		elsif addr = 13 then data <="000000010011";
		elsif addr = 14 then data <="000000010100";
		elsif addr = 15 then data <="000000010101";
		elsif addr = 16 then data <="000000010110";
		elsif addr = 17 then data <="000000010111";
		elsif addr = 18 then data <="000000011000";
		elsif addr = 19 then data <="000000011001";
		elsif addr = 20 then data <="000000100000";
		elsif addr = 21 then data <="000000100001";
		elsif addr = 22 then data <="000000100010";
		elsif addr = 23 then data <="000000100011";
		elsif addr = 24 then data <="000000100100";
		elsif addr = 25 then data <="000000100101";
		elsif addr = 26 then data <="000000100110";
		elsif addr = 27 then data <="000000100111";
		elsif addr = 28 then data <="000000101000";
		elsif addr = 29 then data <="000000101001";
		elsif addr = 30 then data <="000000110000";
		elsif addr = 31 then data <="000000110001";
		elsif addr = 32 then data <="000000110010";
		elsif addr = 33 then data <="000000110011";
		elsif addr = 34 then data <="000000110100";
		elsif addr = 35 then data <="000000110101";
		elsif addr = 36 then data <="000000110110";
		elsif addr = 37 then data <="000000110111";
		elsif addr = 38 then data <="000000111000";
		elsif addr = 39 then data <="000000111001";
		elsif addr = 40 then data <="000001000000";
		elsif addr = 41 then data <="000001000001";
		elsif addr = 42 then data <="000001000010";
		elsif addr = 43 then data <="000001000011";
		elsif addr = 44 then data <="000001000100";
		elsif addr = 45 then data <="000001000101";
		elsif addr = 46 then data <="000001000110";
		elsif addr = 47 then data <="000001000111";
		elsif addr = 48 then data <="000001001000";
		elsif addr = 49 then data <="000001001001";
		elsif addr = 50 then data <="000001010000";
		elsif addr = 51 then data <="000001010001";
		elsif addr = 52 then data <="000001010010";
		elsif addr = 53 then data <="000001010011";
		elsif addr = 54 then data <="000001010100";
		elsif addr = 55 then data <="000001010101";
		elsif addr = 56 then data <="000001010110";
		elsif addr = 57 then data <="000001010111";
		elsif addr = 58 then data <="000001011000";
		elsif addr = 59 then data <="000001011001";
		elsif addr = 60 then data <="000001100000";
		elsif addr = 61 then data <="000001100001";
		elsif addr = 62 then data <="000001100010";
		elsif addr = 63 then data <="000001100011";
		elsif addr = 64 then data <="000001100100";
		elsif addr = 65 then data <="000001100101";
		elsif addr = 66 then data <="000001100110";
		elsif addr = 67 then data <="000001100111";
		elsif addr = 68 then data <="000001101000";
		elsif addr = 69 then data <="000001101001";
		elsif addr = 70 then data <="000001110000";
		elsif addr = 71 then data <="000001110001";
		elsif addr = 72 then data <="000001110010";
		elsif addr = 73 then data <="000001110011";
		elsif addr = 74 then data <="000001110100";
		elsif addr = 75 then data <="000001110101";
		elsif addr = 76 then data <="000001110110";
		elsif addr = 77 then data <="000001110111";
		elsif addr = 78 then data <="000001111000";
		elsif addr = 79 then data <="000001111001";
		elsif addr = 80 then data <="000010000000";
		elsif addr = 81 then data <="000010000001";
		elsif addr = 82 then data <="000010000010";
		elsif addr = 83 then data <="000010000011";
		elsif addr = 84 then data <="000010000100";
		elsif addr = 85 then data <="000010000101";
		elsif addr = 86 then data <="000010000110";
		elsif addr = 87 then data <="000010000111";
		elsif addr = 88 then data <="000010001000";
		elsif addr = 89 then data <="000010001001";
		elsif addr = 90 then data <="000010010000";
		elsif addr = 91 then data <="000010010001";
		elsif addr = 92 then data <="000010010010";
		elsif addr = 93 then data <="000010010011";
		elsif addr = 94 then data <="000010010100";
		elsif addr = 95 then data <="000010010101";
		elsif addr = 96 then data <="000010010110";
		elsif addr = 97 then data <="000010010111";
		elsif addr = 98 then data <="000010011000";
		elsif addr = 99 then data <="000010011001";
		elsif addr = 100 then data <="000000000000";
		elsif addr = 101 then data <="000100000001";
		elsif addr = 102 then data <="000100000010";
		elsif addr = 103 then data <="000100000011";
		elsif addr = 104 then data <="000100000100";
		elsif addr = 105 then data <="000100000101";
		elsif addr = 106 then data <="000100000110";
		elsif addr = 107 then data <="000100000111";
		elsif addr = 108 then data <="000100001000";
		elsif addr = 109 then data <="000100001001";
		elsif addr = 110 then data <="000100010000";
		elsif addr = 111 then data <="000100010001";
		elsif addr = 112 then data <="000100010010";
		elsif addr = 113 then data <="000100010011";
		elsif addr = 114 then data <="000100010100";
		elsif addr = 115 then data <="000100010101";
		elsif addr = 116 then data <="000100010110";
		elsif addr = 117 then data <="000100010111";
		elsif addr = 118 then data <="000100011000";
		elsif addr = 119 then data <="000100011001";
		elsif addr = 120 then data <="000100100000";
		elsif addr = 121 then data <="000100100001";
		elsif addr = 122 then data <="000100100010";
		elsif addr = 123 then data <="000100100011";
		elsif addr = 124 then data <="000100100100";
		elsif addr = 125 then data <="000100100101";
		elsif addr = 126 then data <="000100100110";
		elsif addr = 127 then data <="000100100111";
		elsif addr = 128 then data <="000100101000";
		elsif addr = 129 then data <="000100101001";
		elsif addr = 130 then data <="000100110000";
		elsif addr = 131 then data <="000100110001";
		elsif addr = 132 then data <="000100110010";
		elsif addr = 133 then data <="000100110011";
		elsif addr = 134 then data <="000100110100";
		elsif addr = 135 then data <="000100110101";
		elsif addr = 136 then data <="000100110110";
		elsif addr = 137 then data <="000100110111";
		elsif addr = 138 then data <="000100111000";
		elsif addr = 139 then data <="000100111001";
		elsif addr = 140 then data <="000101000000";
		elsif addr = 141 then data <="000101000001";
		elsif addr = 142 then data <="000101000010";
		elsif addr = 143 then data <="000101000011";
		elsif addr = 144 then data <="000101000100";
		elsif addr = 145 then data <="000101000101";
		elsif addr = 146 then data <="000101000110";
		elsif addr = 147 then data <="000101000111";
		elsif addr = 148 then data <="000101001000";
		elsif addr = 149 then data <="000101001001";
		elsif addr = 150 then data <="000101010000";
		elsif addr = 151 then data <="000101010001";
		elsif addr = 152 then data <="000101010010";
		elsif addr = 153 then data <="000101010011";
		elsif addr = 154 then data <="000101010100";
		elsif addr = 155 then data <="000101010101";
		elsif addr = 156 then data <="000101010110";
		elsif addr = 157 then data <="000101010111";
		elsif addr = 158 then data <="000101011000";
		elsif addr = 159 then data <="000101011001";
		elsif addr = 160 then data <="000101100000";
		elsif addr = 161 then data <="000101100001";
		elsif addr = 162 then data <="000101100010";
		elsif addr = 163 then data <="000101100011";
		elsif addr = 164 then data <="000101100100";
		elsif addr = 165 then data <="000101100101";
		elsif addr = 166 then data <="000101100110";
		elsif addr = 167 then data <="000101100111";
		elsif addr = 168 then data <="000101101000";
		elsif addr = 169 then data <="000101101001";
		elsif addr = 170 then data <="000101110000";
		elsif addr = 171 then data <="000101110001";
		elsif addr = 172 then data <="000101110010";
		elsif addr = 173 then data <="000101110011";
		elsif addr = 174 then data <="000101110100";
		elsif addr = 175 then data <="000101110101";
		elsif addr = 176 then data <="000101110110";
		elsif addr = 177 then data <="000101110111";
		elsif addr = 178 then data <="000101111000";
		elsif addr = 179 then data <="000101111001";
		elsif addr = 180 then data <="000110000000";
		elsif addr = 181 then data <="000110000001";
		elsif addr = 182 then data <="000110000010";
		elsif addr = 183 then data <="000110000011";
		elsif addr = 184 then data <="000110000100";
		elsif addr = 185 then data <="000110000101";
		elsif addr = 186 then data <="000110000110";
		elsif addr = 187 then data <="000110000111";
		elsif addr = 188 then data <="000110001000";
		elsif addr = 189 then data <="000110001001";
		elsif addr = 190 then data <="000110010000";
		elsif addr = 191 then data <="000110010001";
		elsif addr = 192 then data <="000110010010";
		elsif addr = 193 then data <="000110010011";
		elsif addr = 194 then data <="000110010100";
		elsif addr = 195 then data <="000110010101";
		elsif addr = 196 then data <="000110010110";
		elsif addr = 197 then data <="000110010111";
		elsif addr = 198 then data <="000110011000";
		elsif addr = 199 then data <="000110011001";
		elsif addr = 200 then data <="000100000000";
		elsif addr = 201 then data <="001000000001";
		elsif addr = 202 then data <="001000000010";
		elsif addr = 203 then data <="001000000011";
		elsif addr = 204 then data <="001000000100";
		elsif addr = 205 then data <="001000000101";
		elsif addr = 206 then data <="001000000110";
		elsif addr = 207 then data <="001000000111";
		elsif addr = 208 then data <="001000001000";
		elsif addr = 209 then data <="001000001001";
		elsif addr = 210 then data <="001000010000";
		elsif addr = 211 then data <="001000010001";
		elsif addr = 212 then data <="001000010010";
		elsif addr = 213 then data <="001000010011";
		elsif addr = 214 then data <="001000010100";
		elsif addr = 215 then data <="001000010101";
		elsif addr = 216 then data <="001000010110";
		elsif addr = 217 then data <="001000010111";
		elsif addr = 218 then data <="001000011000";
		elsif addr = 219 then data <="001000011001";
		elsif addr = 220 then data <="001000100000";
		elsif addr = 221 then data <="001000100001";
		elsif addr = 222 then data <="001000100010";
		elsif addr = 223 then data <="001000100011";
		elsif addr = 224 then data <="001000100100";
		elsif addr = 225 then data <="001000100101";
		elsif addr = 226 then data <="001000100110";
		elsif addr = 227 then data <="001000100111";
		elsif addr = 228 then data <="001000101000";
		elsif addr = 229 then data <="001000101001";
		elsif addr = 230 then data <="001000110000";
		elsif addr = 231 then data <="001000110001";
		elsif addr = 232 then data <="001000110010";
		elsif addr = 233 then data <="001000110011";
		elsif addr = 234 then data <="001000110100";
		elsif addr = 235 then data <="001000110101";
		elsif addr = 236 then data <="001000110110";
		elsif addr = 237 then data <="001000110111";
		elsif addr = 238 then data <="001000111000";
		elsif addr = 239 then data <="001000111001";
		elsif addr = 240 then data <="001001000000";
		elsif addr = 241 then data <="001001000001";
		elsif addr = 242 then data <="001001000010";
		elsif addr = 243 then data <="001001000011";
		elsif addr = 244 then data <="001001000100";
		elsif addr = 245 then data <="001001000101";
		elsif addr = 246 then data <="001001000110";
		elsif addr = 247 then data <="001001000111";
		elsif addr = 248 then data <="001001001000";
		elsif addr = 249 then data <="001001001001";
		elsif addr = 250 then data <="001001010000";
		elsif addr = 251 then data <="001001010001";
		elsif addr = 252 then data <="001001010010";
		elsif addr = 253 then data <="001001010011";
		elsif addr = 254 then data <="001001010100";
		elsif addr = 255 then data <="001001010101";
		else data <= "000000000000";
		end if;
	end process;
end behavioural;